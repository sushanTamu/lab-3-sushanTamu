///////////////////////////////////////////////////////////////////////////
// Texas A&M University
// CSCE 616 Hardware Design Verification
// File name   : htax_defines.sv
// Created by  : Prof. Quinn and Saumil Gogri
///////////////////////////////////////////////////////////////////////////


`define PORTS 		4 // Total number of ports in our design are 4
`define VC 				2	// Available virtual channels per port
`define WIDTH			64 //Width on one data packet
